/media/psf/Data/Code/Spectrometer/firmware/speadp/speadp.srcs/sources_1/new/running_generator.vhd